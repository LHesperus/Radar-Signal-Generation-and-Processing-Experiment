library verilog;
use verilog.vl_types.all;
entity altlvds_tx is
    generic(
        number_of_channels: integer := 1;
        deserialization_factor: integer := 4;
        registered_input: string  := "ON";
        multi_clock     : string  := "OFF";
        inclock_period  : integer := 10000;
        outclock_divide_by: vl_notype;
        inclock_boost   : vl_notype;
        center_align_msb: string  := "OFF";
        intended_device_family: string  := "Stratix";
        output_data_rate: integer := 0;
        inclock_data_alignment: string  := "EDGE_ALIGNED";
        outclock_alignment: string  := "EDGE_ALIGNED";
        common_rx_tx_pll: string  := "ON";
        outclock_resource: string  := "AUTO";
        use_external_pll: string  := "OFF";
        implement_in_les: string  := "OFF";
        preemphasis_setting: integer := 0;
        vod_setting     : integer := 0;
        differential_drive: integer := 0;
        outclock_multiply_by: integer := 1;
        coreclock_divide_by: integer := 2;
        outclock_duty_cycle: integer := 50;
        inclock_phase_shift: integer := 0;
        outclock_phase_shift: integer := 0;
        use_no_phase_shift: string  := "ON";
        pll_self_reset_on_loss_lock: string  := "OFF";
        refclk_frequency: string  := "UNUSED";
        data_rate       : string  := "UNUSED";
        lpm_type        : string  := "altlvds_tx";
        lpm_hint        : string  := "UNUSED";
        clk_src_is_pll  : string  := "off";
        STRATIX_TX_STYLE: vl_notype;
        STRATIXII_TX_STYLE: vl_notype;
        CYCLONE_TX_STYLE: vl_notype;
        CYCLONEII_TX_STYLE: vl_notype;
        STRATIXIII_TX_STYLE: vl_notype;
        CYCLONEIII_TX_STYLE: vl_notype;
        MAXV_TX_STYLE   : vl_notype;
        FAMILY_HAS_FLEXIBLE_LVDS: vl_notype;
        FAMILY_HAS_STRATIX_STYLE_PLL: vl_notype;
        FAMILY_HAS_STRATIXII_STYLE_PLL: vl_notype;
        FAMILY_HAS_STRATIXIII_STYLE_PLL: vl_notype;
        INT_CLOCK_BOOST : vl_notype;
        PLL_M_VALUE     : vl_notype;
        PLL_D_VALUE     : vl_notype;
        STRATIX_INCLOCK_BOOST: vl_notype;
        PHASE_INCLOCK   : vl_notype;
        STXII_PHASE_INCLOCK: vl_notype;
        PHASE_OUTCLOCK  : vl_notype;
        STX_PHASE_OUTCLOCK: vl_notype;
        STXII_PHASE_OUTCLOCK: vl_notype;
        STXII_LE_PHASE_INCLOCK: vl_notype;
        STXII_LE_PHASE_OUTCLOCK: vl_notype;
        STXIII_LE_PHASE_INCLOCK: vl_notype;
        STXIII_LE_PHASE_OUTCLOCK: vl_notype;
        REGISTER_WIDTH  : vl_notype;
        FAST_CLK_ENA_PHASE_SHIFT: vl_notype;
        CLOCK_PERIOD    : vl_notype;
        USE_NEW_CORECLK_CKT: vl_notype
    );
    port(
        tx_in           : in     vl_logic_vector;
        tx_inclock      : in     vl_logic;
        tx_syncclock    : in     vl_logic;
        tx_enable       : in     vl_logic;
        sync_inclock    : in     vl_logic;
        tx_pll_enable   : in     vl_logic;
        pll_areset      : in     vl_logic;
        tx_data_reset   : in     vl_logic;
        tx_out          : out    vl_logic_vector;
        tx_outclock     : out    vl_logic;
        tx_coreclock    : out    vl_logic;
        tx_locked       : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of number_of_channels : constant is 1;
    attribute mti_svvh_generic_type of deserialization_factor : constant is 1;
    attribute mti_svvh_generic_type of registered_input : constant is 1;
    attribute mti_svvh_generic_type of multi_clock : constant is 1;
    attribute mti_svvh_generic_type of inclock_period : constant is 1;
    attribute mti_svvh_generic_type of outclock_divide_by : constant is 3;
    attribute mti_svvh_generic_type of inclock_boost : constant is 3;
    attribute mti_svvh_generic_type of center_align_msb : constant is 1;
    attribute mti_svvh_generic_type of intended_device_family : constant is 1;
    attribute mti_svvh_generic_type of output_data_rate : constant is 1;
    attribute mti_svvh_generic_type of inclock_data_alignment : constant is 1;
    attribute mti_svvh_generic_type of outclock_alignment : constant is 1;
    attribute mti_svvh_generic_type of common_rx_tx_pll : constant is 1;
    attribute mti_svvh_generic_type of outclock_resource : constant is 1;
    attribute mti_svvh_generic_type of use_external_pll : constant is 1;
    attribute mti_svvh_generic_type of implement_in_les : constant is 1;
    attribute mti_svvh_generic_type of preemphasis_setting : constant is 1;
    attribute mti_svvh_generic_type of vod_setting : constant is 1;
    attribute mti_svvh_generic_type of differential_drive : constant is 1;
    attribute mti_svvh_generic_type of outclock_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of coreclock_divide_by : constant is 1;
    attribute mti_svvh_generic_type of outclock_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of inclock_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of outclock_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of use_no_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of pll_self_reset_on_loss_lock : constant is 1;
    attribute mti_svvh_generic_type of refclk_frequency : constant is 1;
    attribute mti_svvh_generic_type of data_rate : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of lpm_hint : constant is 1;
    attribute mti_svvh_generic_type of clk_src_is_pll : constant is 1;
    attribute mti_svvh_generic_type of STRATIX_TX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of STRATIXII_TX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of CYCLONE_TX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of CYCLONEII_TX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of STRATIXIII_TX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of CYCLONEIII_TX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of MAXV_TX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of FAMILY_HAS_FLEXIBLE_LVDS : constant is 3;
    attribute mti_svvh_generic_type of FAMILY_HAS_STRATIX_STYLE_PLL : constant is 3;
    attribute mti_svvh_generic_type of FAMILY_HAS_STRATIXII_STYLE_PLL : constant is 3;
    attribute mti_svvh_generic_type of FAMILY_HAS_STRATIXIII_STYLE_PLL : constant is 3;
    attribute mti_svvh_generic_type of INT_CLOCK_BOOST : constant is 3;
    attribute mti_svvh_generic_type of PLL_M_VALUE : constant is 3;
    attribute mti_svvh_generic_type of PLL_D_VALUE : constant is 3;
    attribute mti_svvh_generic_type of STRATIX_INCLOCK_BOOST : constant is 3;
    attribute mti_svvh_generic_type of PHASE_INCLOCK : constant is 3;
    attribute mti_svvh_generic_type of STXII_PHASE_INCLOCK : constant is 3;
    attribute mti_svvh_generic_type of PHASE_OUTCLOCK : constant is 3;
    attribute mti_svvh_generic_type of STX_PHASE_OUTCLOCK : constant is 3;
    attribute mti_svvh_generic_type of STXII_PHASE_OUTCLOCK : constant is 3;
    attribute mti_svvh_generic_type of STXII_LE_PHASE_INCLOCK : constant is 3;
    attribute mti_svvh_generic_type of STXII_LE_PHASE_OUTCLOCK : constant is 3;
    attribute mti_svvh_generic_type of STXIII_LE_PHASE_INCLOCK : constant is 3;
    attribute mti_svvh_generic_type of STXIII_LE_PHASE_OUTCLOCK : constant is 3;
    attribute mti_svvh_generic_type of REGISTER_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of FAST_CLK_ENA_PHASE_SHIFT : constant is 3;
    attribute mti_svvh_generic_type of CLOCK_PERIOD : constant is 3;
    attribute mti_svvh_generic_type of USE_NEW_CORECLK_CKT : constant is 3;
end altlvds_tx;
