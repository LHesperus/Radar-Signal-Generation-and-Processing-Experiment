library verilog;
use verilog.vl_types.all;
entity experiment_tb is
end experiment_tb;
