library verilog;
use verilog.vl_types.all;
entity fir_tb is
end fir_tb;
